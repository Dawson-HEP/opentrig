module clk_ref (
    input wire sampling_clk,

    input wire clk_in_async,
    input wire ref_reset_async,

    output reg [63:0] ref
);
    sync sync_clk_in (
        .async(clk_in_async),
        .clk(sampling_clk),
        .rising(clk_in_rising)
    );
    sync sync_ref_reset (
        .async(ref_reset_async),
        .clk(sampling_clk),
        .falling(ref_reset_falling)
    );

    reg [31:0] low, high;
    reg incr_high;

    always @(posedge sampling_clk) begin
        if (ref_reset_falling) begin
            low <= 0;
            high <= 0;
            incr_high <= 0;
        end else begin
            if (clk_in_rising) begin
                ref <= {high, low};

                if (low == 32'hFFFF_FFFF) begin
                    incr_high <= 1;
                end
                low <= low + 1;
            end else if (incr_high) begin
                high <= high + 1;
                incr_high <= 0;
            end
        end
    end
endmodule
