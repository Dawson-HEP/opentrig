// module trigger_id_parser(
//     input wire 
// );


// endmodule